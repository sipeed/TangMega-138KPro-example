parameter M=32;
parameter N=32;
parameter Q=3;
parameter LATENCY=2;
