`define module_name Ten_Giga_Serial_Ethernet_Top
`define REFCLK0
`define DBG_O
