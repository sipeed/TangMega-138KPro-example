`define Q1_LN0
`define Q1_LN0_PMA_WIDTH 20
`define Q1_LN0_TX_GEARBOX 4
`define Q1_LN0_RX_GEARBOX 4
`define Q1_LN0_8B10B_ENCODE
`define Q1_LN0_8B10B_DECODE
`define Q1_LN0_WORD_ALIGN
`define Q1_LN0_CHANNEL_BONDING_MASTER_SEL 0
`define Q1_LN0_TX_IF_MST_SEL 0
`define Q1_LN1
`define Q1_LN1_PMA_WIDTH 20
`define Q1_LN1_TX_GEARBOX 4
`define Q1_LN1_RX_GEARBOX 4
`define Q1_LN1_8B10B_ENCODE
`define Q1_LN1_8B10B_DECODE
`define Q1_LN1_WORD_ALIGN
`define Q1_LN1_CHANNEL_BONDING_MASTER_SEL 0
`define Q1_LN1_TX_IF_MST_SEL 0
`define MODULE_NAME Customized_PHY_Top
