`define module_name Ten_Giga_Serial_Ethernet_Top_1
`define REFCLK0
`define DBG_O
